LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DISPLAY IS
    PORT(M:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    BCD:OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
    END DISPLAY;
ARCHITECTURE A OF DISPLAY IS
    BEGIN
PROCESS(M)
BEGIN
    CASE M IS
    WHEN "0000"=>BCD<="1000000";
    WHEN "0001"=>BCD<="1111001";
    WHEN "0010"=>BCD<="0100100";
    WHEN "0011"=>BCD<="0110000";
    WHEN "0100"=>BCD<="0011001";
    WHEN "0101"=>BCD<="0010010";
    WHEN "0110"=>BCD<="0000010";
    WHEN "0111"=>BCD<="1111000";
    WHEN "1000"=>BCD<="0000000";
    WHEN "1001"=>BCD<="0010000";
WHEN OTHERS => BCD <="1111111";
END CASE;
END PROCESS;
END A;
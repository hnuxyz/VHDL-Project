LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY FASHENG IS
PORT(CLK1,CLR,EN:IN STD_LOGIC;
    SOUND:OUT STD_LOGIC);
END FASHENG;
ARCHITECTURE A OF FASHENG IS
    BEGIN
PROCESS(EN,CLK1)
BEGIN
IF(CLK1'EVENT AND CLK1='1') THEN
    IF(CLR='0' AND EN='1') THEN
        SOUND<='1';
    ELSE
        SOUND<='0';
    END IF;
END IF;
END PROCESS;
END A;
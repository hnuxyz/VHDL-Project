LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY FENPIN IS
	PORT(CLK:IN STD_LOGIC;
		CLK1:OUT STD_LOGIC);
END FENPIN;
ARCHITECTURE clk_div_behavior OF FENPIN IS
	SIGNAL counter:STD_LOGIC_VECTOR(24 DOWNTO 0);
	SIGNAL temp:STD_LOGIC;
BEGIN
	PROCESS(CLK)
	BEGIN
		IF(CLK'EVENT AND CLK='1')THEN
			IF(counter="1011111010111100000111111")THEN       
				counter<="0000000000000000000000000";
				temp<=NOT temp;
			ELSE
				counter<=counter+1;
			END	IF;
		END IF;
	END PROCESS;
	CLK1<=temp;
END clk_div_behavior;



LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DJSQ IS
PORT(CLR,CLK1,EN:IN STD_LOGIC;
	H,L:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	SOUND1:OUT STD_LOGIC);
END DJSQ;
ARCHITECTURE DJSQ_ARC OF DJSQ IS
BEGIN
PROCESS(CLK1,EN)
VARIABLE HH,LL:STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
IF CLR='0' THEN
HH:="0011";
LL:="0000";
ELSE
IF CLK1'EVENT AND CLK1='1'THEN
IF EN='0'THEN
IF LL=0 AND HH=0 THEN
SOUND1<='1';
ELSIF LL=0 THEN
LL:="1001";
HH:=HH-1;
ELSE
LL:=LL-1;
END IF;
ELSE
SOUND1<='0';
HH:="0011";
LL:="0000";
END IF;
END IF;
END IF;
H<=HH;
L<=LL;
END PROCESS;
END DJSQ_ARC;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DISPLAY1 IS
    PORT(H,L:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    BCD1,BCD2:OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
    END DISPLAY1;
ARCHITECTURE B OF DISPLAY1 IS
    BEGIN
PROCESS(H)
BEGIN
    CASE H IS
    WHEN "0000"=>BCD1<="1000000";
    WHEN "0001"=>BCD1<="1111001";
    WHEN "0010"=>BCD1<="0100100";
    WHEN "0011"=>BCD1<="0110000";
    WHEN "0100"=>BCD1<="0011001";
    WHEN "0101"=>BCD1<="0010010";
    WHEN "0110"=>BCD1<="0000010";
    WHEN "0111"=>BCD1<="1111000";
    WHEN "1000"=>BCD1<="0000000";
    WHEN "1001"=>BCD1<="0010000";
WHEN OTHERS => BCD1 <="1111111";
END CASE;
END PROCESS;
PROCESS(L)
BEGIN
    CASE L IS
    WHEN "0000"=>BCD2<="1000000";
    WHEN "0001"=>BCD2<="1111001";
    WHEN "0010"=>BCD2<="0100100";
    WHEN "0011"=>BCD2<="0110000";
    WHEN "0100"=>BCD2<="0011001";
    WHEN "0101"=>BCD2<="0010010";
    WHEN "0110"=>BCD2<="0000010";
    WHEN "0111"=>BCD2<="1111000";
    WHEN "1000"=>BCD2<="0000000";
    WHEN "1001"=>BCD2<="0010000";
WHEN OTHERS => BCD2 <="1111111";
END CASE;
END PROCESS;
END B;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY QDJB IS
PORT(S1,S2,S3,S4,S5,S6,S7,S8,CLR,OE:IN STD_LOGIC;
	  Q1,Q2,Q3,Q4,Q5,Q6,Q7,Q8:OUT STD_LOGIC);
END QDJB;
ARCHITECTURE A OF QDJB IS
	BEGIN
PROCESS(S1,S2,S3,S4,S5,S6,S7,S8,OE,CLR)
BEGIN
IF(CLR='1')THEN
Q1<='0';Q2<='0';Q3<='0';Q4<='0';Q5<='0';Q6<='0';Q7<='0';Q8<='0';
ELSIF(OE='0')THEN
Q1<=S1;Q2<=S2;Q3<=S3;Q4<=S4;Q5<=S5;Q6<=S6;Q7<=S7;Q8<=S8;
END IF;
END PROCESS;
END A;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY BIANMA IS
PORT(Q1,Q2,Q3,Q4,Q5,Q6,Q7,Q8:IN STD_LOGIC;
	CLR:IN STD_LOGIC;
	M:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	EN:OUT STD_LOGIC);
END BIANMA;
ARCHITECTURE A OF BIANMA IS
BEGIN
PROCESS(Q1,Q2,Q3,Q4,Q5,Q6,Q7,Q8,CLR)
VARIABLE TEMP: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
TEMP:=Q1&Q2&Q3&Q4&Q5&Q6&Q7&Q8;
CASE TEMP IS
WHEN"10000000"=>M<="0001";
WHEN"01000000"=>M<="0010";
WHEN"00100000"=>M<="0011";
WHEN"00010000"=>M<="0100";
WHEN"00001000"=>M<="0101";
WHEN"00000100"=>M<="0110";
WHEN"00000010"=>M<="0111";
WHEN"00000001"=>M<="1000";
WHEN OTHERS=>M<="1111";
END CASE;
EN <=TEMP(7) OR TEMP(6) OR TEMP(5) OR TEMP(4) OR TEMP(3) OR TEMP(2) OR TEMP(1) OR TEMP(0) OR CLR;
END PROCESS;
END A; 